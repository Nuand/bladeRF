-- Copyright (c) 2013 Nuand LLC
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
-- THE SOFTWARE.

library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.math_real.all;
    use ieee.math_complex.all;

library work;
    use work.bladerf_p.all;

architecture hosted_bladerf of bladerf is

    attribute noprune          : boolean;
    attribute keep             : boolean;

    alias  sys_reset_async     : std_logic is fx3_ctl(7);
    signal sys_reset_pclk      : std_logic;
    signal sys_reset           : std_logic;

    signal sys_clock           : std_logic;
    signal sys_pll_locked      : std_logic;
    signal sys_pll_reset       : std_logic;

    signal fx3_pclk_pll        : std_logic;
    signal fx3_pclk_pll_locked : std_logic;
    signal fx3_pclk_pll_reset  : std_logic;

    -- Can be set from libbladeRF using bladerf_set_rx_mux()
    type rx_mux_mode_t is (
        RX_MUX_NORMAL,
        RX_MUX_12BIT_COUNTER,
        RX_MUX_32BIT_COUNTER,
        RX_MUX_ENTROPY,
        RX_MUX_DIGITAL_LOOPBACK
    );

    signal rx_mux_mode           : rx_mux_mode_t;
    signal rx_mux_sel            : unsigned(2 downto 0);

    signal nios_gpio_i           : std_logic_vector(31 downto 0);
    signal nios_xb_gpio_in       : std_logic_vector(31 downto 0) := (others => '0');
    signal nios_xb_gpio_out      : std_logic_vector(31 downto 0) := (others => '0');
    signal nios_xb_gpio_oe       : std_logic_vector(31 downto 0) := (others => '0');

    signal nios_gpio             : nios_gpio_t;

    signal i2c_scl_in            : std_logic;
    signal i2c_scl_out           : std_logic;
    signal i2c_scl_oen           : std_logic;

    signal i2c_sda_in            : std_logic;
    signal i2c_sda_out           : std_logic;
    signal i2c_sda_oen           : std_logic;

    signal rx_sample_fifo        : fifo_t := FIFO_T_DEFAULT;
    signal tx_sample_fifo        : fifo_t := FIFO_T_DEFAULT;
    signal rx_loopback_fifo      : fifo_t := FIFO_T_DEFAULT;

    signal tx_meta_fifo          : meta_fifo_tx_t := META_FIFO_TX_T_DEFAULT;
    signal rx_meta_fifo          : meta_fifo_rx_t := META_FIFO_RX_T_DEFAULT;

    signal usb_speed_pclk        : std_logic;
    signal usb_speed_rx          : std_logic;
    signal usb_speed_tx          : std_logic;

    signal tx_reset              : std_logic;
    signal rx_reset              : std_logic;

    signal tx_enable_pclk        : std_logic;
    signal rx_enable_pclk        : std_logic;

    signal tx_enable             : std_logic;
    signal rx_enable             : std_logic;

    signal meta_en_tx            : std_logic;
    signal meta_en_rx            : std_logic;
    signal meta_en_pclk          : std_logic;

    signal tx_timestamp          : unsigned(63 downto 0);
    signal rx_timestamp          : unsigned(63 downto 0);
    signal timestamp_sync        : std_logic;

    signal rx_sample_i           : signed(15 downto 0);
    signal rx_sample_q           : signed(15 downto 0);
    signal rx_sample_valid       : std_logic;

    signal rx_gen_mode           : std_logic;
    signal rx_gen_i              : signed(15 downto 0);
    signal rx_gen_q              : signed(15 downto 0);
    signal rx_gen_valid          : std_logic;

    signal rx_loopback_i         : signed(15 downto 0) := (others =>'0');
    signal rx_loopback_q         : signed(15 downto 0) := (others =>'0');
    signal rx_loopback_valid     : std_logic := '0';
    signal rx_loopback_enabled   : std_logic := '0';
    signal tx_loopback_enabled   : std_logic := '0';

    signal tx_sample_i           : signed(15 downto 0);
    signal tx_sample_q           : signed(15 downto 0);
    signal tx_sample_valid       : std_logic;

    signal fx3_gpif_in           : std_logic_vector(31 downto 0);
    signal fx3_gpif_out          : std_logic_vector(31 downto 0);
    signal fx3_gpif_oe           : std_logic;

    signal fx3_ctl_in            : std_logic_vector(12 downto 0);
    signal fx3_ctl_out           : std_logic_vector(12 downto 0);
    signal fx3_ctl_oe            : std_logic_vector(12 downto 0);

    signal tx_underflow_led      : std_logic := '1';

    signal rx_overflow_led       : std_logic := '1';

    signal rx_mux_i              : signed(15 downto 0);
    signal rx_mux_q              : signed(15 downto 0);
    signal rx_mux_valid          : std_logic;

    signal led1_blink            : std_logic;

    signal nios_sdo              : std_logic;
    signal nios_sdio             : std_logic;
    signal nios_sclk             : std_logic;
    signal nios_ss_n             : std_logic_vector(1 downto 0);

    signal command_serial_in     : std_logic;
    signal command_serial_out    : std_logic;

    signal timestamp_req         : std_logic;
    signal timestamp_ack         : std_logic;
    signal fx3_timestamp         : unsigned(63 downto 0);

    signal rx_ts_reset           : std_logic;
    signal tx_ts_reset           : std_logic;

    -- Trigger Control interfaces
    signal rx_trigger_ctl        : std_logic_vector(7 downto 0);
    signal tx_trigger_ctl        : std_logic_vector(7 downto 0);

    -- Trigger Control breakdown
    alias rx_trigger_arm         : std_logic is rx_trigger_ctl(0);
    alias rx_trigger_fire        : std_logic is rx_trigger_ctl(1);
    alias rx_trigger_master      : std_logic is rx_trigger_ctl(2);
    alias rx_trigger_line        : std_logic is mini_exp1;
    signal rx_trigger_signal_out : std_logic := '0';

    alias tx_trigger_arm         : std_logic is tx_trigger_ctl(0);
    alias tx_trigger_fire        : std_logic is tx_trigger_ctl(1);
    alias tx_trigger_master      : std_logic is tx_trigger_ctl(2);
    alias tx_trigger_line        : std_logic is mini_exp1;

    signal tx_trigger_arm_sync   : std_logic;
    signal tx_trigger_line_sync  : std_logic;

    -- Trigger Control readback interfaces
    signal rx_trigger_ctl_rb     : std_logic_vector(7 downto 0);
    signal tx_trigger_ctl_rb     : std_logic_vector(7 downto 0);

    -- Trigger Control readback breakdown
    alias rx_trigger_arm_rb      : std_logic is rx_trigger_ctl_rb(0);
    alias rx_trigger_fire_rb     : std_logic is rx_trigger_ctl_rb(1);
    alias rx_trigger_master_rb   : std_logic is rx_trigger_ctl_rb(2);
    alias rx_trigger_line_rb     : std_logic is rx_trigger_ctl_rb(3);
    alias rx_trigger_unused_rb   : std_logic_vector(7 downto 4) is rx_trigger_ctl_rb(7 downto 4);

    alias tx_trigger_arm_rb      : std_logic is tx_trigger_ctl_rb(0);
    alias tx_trigger_fire_rb     : std_logic is tx_trigger_ctl_rb(1);
    alias tx_trigger_master_rb   : std_logic is tx_trigger_ctl_rb(2);
    alias tx_trigger_line_rb     : std_logic is tx_trigger_ctl_rb(3);
    alias tx_trigger_unused_rb   : std_logic_vector(7 downto 4) is tx_trigger_ctl_rb(7 downto 4);

    -- Trigger Outputs
    signal lms_rx_enable_sig                 : std_logic;
    signal lms_rx_enable_qualified           : std_logic;
    signal tx_sample_fifo_rempty_untriggered : std_logic;

    signal tx_lms_data     : signed(11 downto 0) := (others => '0');

    signal rffe_gpio       : rffe_gpio_t := (
        i => RFFE_GPI_DEFAULT,
        o => pack(RFFE_GPO_DEFAULT)
    );

    signal ad9361 : mimo_2r2t_t := MIMO_2R2T_T_DEFAULT;
    alias tx_clock  is ad9361.clock;
    alias rx_clock  is ad9361.clock;

    signal channel_sel : std_logic := '0';

begin

    -- ========================================================================
    -- PLLs
    -- ========================================================================

    -- Create 80 MHz system clock from c5_clock_1 (38.4 MHz)
    U_system_pll : component system_pll
        port map (
            refclk   => c5_clock_1,
            rst      => sys_pll_reset,
            outclk_0 => sys_clock,
            locked   => sys_pll_locked
        );

    U_pll_reset_pll : entity work.pll_reset
        generic map (
            SYS_CLOCK_FREQ_HZ   => 38_400_000,
            DEVICE_FAMILY       => "Cyclone V"
        )
        port map (
            sys_clock      => c5_clock_1,
            pll_locked     => sys_pll_locked,
            pll_reset      => sys_pll_reset
        );

    -- Use PLL to adjust the phase of the FX3 PCLK to
    -- retime the FX3 GPIF interface for timing closure.
    U_fx3_pll : component fx3_pll
        port map (
            refclk   =>  fx3_pclk,
            rst      =>  fx3_pclk_pll_reset,
            outclk_0 =>  fx3_pclk_pll,
            locked   =>  fx3_pclk_pll_locked
        );

    U_pll_reset_fx3_pll : entity work.pll_reset
        generic map (
            SYS_CLOCK_FREQ_HZ   => 100_000_000,
            DEVICE_FAMILY       => "Cyclone V"
        )
        port map (
            sys_clock      => fx3_pclk,
            pll_locked     => fx3_pclk_pll_locked,
            pll_reset      => fx3_pclk_pll_reset
        );


    -- ========================================================================
    -- POWER SUPPLY SYNCHRONIZATION
    -- ========================================================================

    -- ADP2384 sync freq must be +/- 10% of the Fsw set by RT.
    -- RT = 53.6k +/- 1%, so Fsw = 0.999768 MHz to 1.015514 MHz.
    -- Therefore, sync must fall between:
    --   -10% of 1.015514 MHz = 0.913964 MHz
    --   +10% of 0.999768 MHz = 1.099745 MHz
    -- Dividing 38.4 MHz by 38 yields 1.010526 MHz.
    ps_sync : process(c5_clock_1)
        variable count  : natural range 0 to 19 := 19;
        variable ps_clk : std_logic := '0';
    begin
        if( rising_edge(c5_clock_1) ) then
            ps_sync_1p1 <= ps_clk;
            ps_sync_1p8 <= ps_clk;
            count := count - 1;
            if( count = 0 ) then
                count  := 19;
                ps_clk := not ps_clk;
            end if;
        end if;
    end process;

    -- ========================================================================
    -- FX3 GPIF
    -- ========================================================================

    -- FX3 GPIF
    U_fx3_gpif : entity work.fx3_gpif
        port map (
            pclk                =>  fx3_pclk_pll,
            reset               =>  sys_reset_pclk,

            usb_speed           =>  usb_speed_pclk,

            meta_enable         =>  meta_en_pclk,
            rx_enable           =>  rx_enable_pclk,
            tx_enable           =>  tx_enable_pclk,

            gpif_in             =>  fx3_gpif_in,
            gpif_out            =>  fx3_gpif_out,
            gpif_oe             =>  fx3_gpif_oe,
            ctl_in              =>  fx3_ctl_in,
            ctl_out             =>  fx3_ctl_out,
            ctl_oe              =>  fx3_ctl_oe,

            tx_fifo_write       =>  tx_sample_fifo.wreq,
            tx_fifo_full        =>  tx_sample_fifo.wfull,
            tx_fifo_empty       =>  tx_sample_fifo.wempty,
            tx_fifo_usedw       =>  tx_sample_fifo.wused,
            tx_fifo_data        =>  tx_sample_fifo.wdata,

            tx_timestamp        =>  fx3_timestamp,
            tx_meta_fifo_write  =>  tx_meta_fifo.wreq,
            tx_meta_fifo_full   =>  tx_meta_fifo.wfull,
            tx_meta_fifo_empty  =>  tx_meta_fifo.wempty,
            tx_meta_fifo_usedw  =>  tx_meta_fifo.wused,
            tx_meta_fifo_data   =>  tx_meta_fifo.wdata,

            rx_fifo_read        =>  rx_sample_fifo.rreq,
            rx_fifo_full        =>  rx_sample_fifo.rfull,
            rx_fifo_empty       =>  rx_sample_fifo.rempty,
            rx_fifo_usedw       =>  rx_sample_fifo.rused,
            rx_fifo_data        =>  rx_sample_fifo.rdata,

            rx_meta_fifo_read   =>  rx_meta_fifo.rreq,
            rx_meta_fifo_full   =>  rx_meta_fifo.rfull,
            rx_meta_fifo_empty  =>  rx_meta_fifo.rempty,
            rx_meta_fifo_usedr  =>  rx_meta_fifo.rused,
            rx_meta_fifo_data   =>  rx_meta_fifo.rdata
        );

    -- FX3 GPIF bidirectional signals
    register_gpif : process(sys_reset_pclk, fx3_pclk_pll)
    begin
        if( sys_reset_pclk = '1' ) then
            fx3_gpif    <= (others =>'Z');
            fx3_gpif_in <= (others =>'0');
        elsif( rising_edge(fx3_pclk_pll) ) then
            fx3_gpif_in <= fx3_gpif;
            if( fx3_gpif_oe = '1' ) then
                fx3_gpif <= fx3_gpif_out;
            else
                fx3_gpif <= (others =>'Z');
            end if;
        end if;
    end process;

    -- FX3 CTL bidirectional signals
    generate_ctl : for i in fx3_ctl'range generate
        fx3_ctl(i) <= fx3_ctl_out(i) when fx3_ctl_oe(i) = '1' else 'Z';
    end generate;

    fx3_ctl_in <= fx3_ctl;

    toggle_led1 : process(fx3_pclk_pll)
        variable count : natural range 0 to 10_000_000 := 10_000_000;
    begin
        if( rising_edge(fx3_pclk_pll) ) then
            count := count - 1;
            if( count = 0 ) then
                count := 10_000_000;
                led1_blink <= not led1_blink;
            end if;
        end if;
    end process;


    -- ========================================================================
    -- NIOS SYSTEM
    -- ========================================================================

    U_nios_system : component nios_system
      port map (
        clk_clk                         => sys_clock,
        reset_reset_n                   => '1',
        dac_MISO                        => nios_sdo,
        dac_MOSI                        => nios_sdio,
        dac_SCLK                        => nios_sclk,
        dac_SS_n                        => nios_ss_n,
        spi_MISO                        => adi_spi_sdo,
        spi_MOSI                        => adi_spi_sdi,
        spi_SCLK                        => adi_spi_sclk,
        spi_SS_n                        => adi_spi_csn,
        gpio_export                     => nios_gpio_i,
        gpio_rffe_0_in_port             => pack(rffe_gpio),
        gpio_rffe_0_out_port            => rffe_gpio.o,
        ad9361_dac_sync_in_sync         => '0',
        ad9361_dac_sync_out_sync        => adi_sync_in,
        ad9361_data_clock_clk           => ad9361.clock, -- out std_logic;
        ad9361_data_reset_reset         => ad9361.reset, -- out std_logic;
        ad9361_device_if_rx_clk_in_p    => adi_rx_clock,
        ad9361_device_if_rx_clk_in_n    => '0',
        ad9361_device_if_rx_frame_in_p  => adi_rx_frame,
        ad9361_device_if_rx_frame_in_n  => '0',
        ad9361_device_if_rx_data_in_p   => adi_rx_data,
        ad9361_device_if_rx_data_in_n   => (others => '0'),
        ad9361_device_if_tx_clk_out_p   => adi_tx_clock,
        ad9361_device_if_tx_clk_out_n   => open,
        ad9361_device_if_tx_frame_out_p => adi_tx_frame,
        ad9361_device_if_tx_frame_out_n => open,
        ad9361_device_if_tx_data_out_p  => adi_tx_data,
        ad9361_device_if_tx_data_out_n  => open,
        ad9361_adc_i0_enable            => ad9361.ch(0).adc.i.enable, -- out sl
        ad9361_adc_i0_valid             => ad9361.ch(0).adc.i.valid,  -- out sl
        ad9361_adc_i0_data              => ad9361.ch(0).adc.i.data,   -- out slv(15:0)
        ad9361_adc_i1_enable            => ad9361.ch(1).adc.i.enable, -- out sl
        ad9361_adc_i1_valid             => ad9361.ch(1).adc.i.valid,  -- out sl
        ad9361_adc_i1_data              => ad9361.ch(1).adc.i.data,   -- out slv(15:0)
        ad9361_adc_overflow_ovf         => ad9361.adc_overflow,       -- in  sl
        ad9361_adc_q0_enable            => ad9361.ch(0).adc.q.enable, -- out sl
        ad9361_adc_q0_valid             => ad9361.ch(0).adc.q.valid,  -- out sl
        ad9361_adc_q0_data              => ad9361.ch(0).adc.q.data,   -- out slv(15:0)
        ad9361_adc_q1_enable            => ad9361.ch(1).adc.q.enable, -- out sl
        ad9361_adc_q1_valid             => ad9361.ch(1).adc.q.valid,  -- out sl
        ad9361_adc_q1_data              => ad9361.ch(1).adc.q.data,   -- out slv(15:0)
        ad9361_adc_underflow_unf        => ad9361.adc_underflow,      -- in  sl
        ad9361_dac_i0_enable            => ad9361.ch(0).dac.i.enable, -- out sl
        ad9361_dac_i0_valid             => ad9361.ch(0).dac.i.valid,  -- out sl
        ad9361_dac_i0_data              => ad9361.ch(0).dac.i.data,   -- in  slv(15:0)
        ad9361_dac_i1_enable            => ad9361.ch(1).dac.i.enable, -- out sl
        ad9361_dac_i1_valid             => ad9361.ch(1).dac.i.valid,  -- out sl
        ad9361_dac_i1_data              => ad9361.ch(1).dac.i.data,   -- in  slv(15:0)
        ad9361_dac_overflow_ovf         => ad9361.dac_overflow,       -- in  sl
        ad9361_dac_q0_enable            => ad9361.ch(0).dac.q.enable, -- out sl
        ad9361_dac_q0_valid             => ad9361.ch(0).dac.q.valid,  -- out sl
        ad9361_dac_q0_data              => ad9361.ch(0).dac.q.data,   -- in  slv(15:0)
        ad9361_dac_q1_enable            => ad9361.ch(1).dac.q.enable, -- out sl
        ad9361_dac_q1_valid             => ad9361.ch(1).dac.q.valid,  -- out sl
        ad9361_dac_q1_data              => ad9361.ch(1).dac.q.data,   -- in  slv(15:0)
        ad9361_dac_underflow_unf        => ad9361.dac_underflow,      -- in  sl
        xb_gpio_in_port                 => nios_xb_gpio_in,
        xb_gpio_out_port                => nios_xb_gpio_out,
        xb_gpio_dir_export              => nios_xb_gpio_oe,
        command_serial_in               => command_serial_in,
        command_serial_out              => command_serial_out,
        oc_i2c_arst_i                   => '0',
        oc_i2c_scl_pad_i                => i2c_scl_in,
        oc_i2c_scl_pad_o                => i2c_scl_out,
        oc_i2c_scl_padoen_o             => i2c_scl_oen,
        oc_i2c_sda_pad_i                => i2c_sda_in,
        oc_i2c_sda_pad_o                => i2c_sda_out,
        oc_i2c_sda_padoen_o             => i2c_sda_oen,
        rx_tamer_ts_sync_in             => '0',
        rx_tamer_ts_sync_out            => open,
        rx_tamer_ts_pps                 => '0',
        rx_tamer_ts_clock               => rx_clock,
        rx_tamer_ts_reset               => rx_ts_reset,
        unsigned(rx_tamer_ts_time)      => rx_timestamp,
        tx_tamer_ts_sync_in             => '0',
        tx_tamer_ts_sync_out            => open,
        tx_tamer_ts_pps                 => '0',
        tx_tamer_ts_clock               => tx_clock,
        tx_tamer_ts_reset               => tx_ts_reset,
        unsigned(tx_tamer_ts_time)      => tx_timestamp,
        rx_trigger_ctl_out_port         => rx_trigger_ctl,
        tx_trigger_ctl_out_port         => tx_trigger_ctl,
        rx_trigger_ctl_in_port          => rx_trigger_ctl_rb,
        tx_trigger_ctl_in_port          => tx_trigger_ctl_rb
      );

    -- FX3 UART
    command_serial_in <= fx3_uart_txd       when sys_reset = '0' else '1';
    fx3_uart_rxd      <= command_serial_out when sys_reset = '0' else 'Z';

    -- FX3 UART CTS and Flash SPI CSx are tied to the same signal.
    -- Allow SPI accesses when FPGA is in reset
    fx3_uart_cts      <= '1' when sys_reset_pclk = '0' else 'Z';

    -- Nios GPIO
    nios_gpio.usb_speed   <= nios_gpio_i(7);
    nios_gpio.rx_mux_sel  <= nios_gpio_i(10 downto 8);
    nios_gpio.spi_mux     <= nios_gpio_i(11);
    nios_gpio.leds        <= nios_gpio_i(14 downto 12);
    nios_gpio.led_mode    <= nios_gpio_i(15);
    nios_gpio.meta_sync   <= nios_gpio_i(16);
    nios_gpio.channel_sel <= nios_gpio_i(17);
    nios_gpio.xb_mode     <= nios_gpio_i(31 downto 30);

    -- RFFE GPIO outputs
    adi_ctrl_in    <= unpack(rffe_gpio.o).ctrl_in;
    adi_tx_spdt2_v <= unpack(rffe_gpio.o).tx_spdt2;
    adi_tx_spdt1_v <= unpack(rffe_gpio.o).tx_spdt1;
    tx_bias_en     <= unpack(rffe_gpio.o).tx_bias_en;
    adi_rx_spdt2_v <= unpack(rffe_gpio.o).rx_spdt2;
    adi_rx_spdt1_v <= unpack(rffe_gpio.o).rx_spdt1;
    rx_bias_en     <= unpack(rffe_gpio.o).rx_bias_en;
    --adi_sync_in    <= unpack(rffe_gpio.o).sync_in;
    adi_en_agc     <= unpack(rffe_gpio.o).en_agc;
    adi_txnrx      <= unpack(rffe_gpio.o).txnrx;
    adi_enable     <= unpack(rffe_gpio.o).enable;
    adi_reset_n    <= unpack(rffe_gpio.o).reset_n;

    -- LEDs
    led(1) <= led1_blink        when nios_gpio.led_mode = '0' else not nios_gpio.leds(1);
    led(2) <= tx_underflow_led  when nios_gpio.led_mode = '0' else not nios_gpio.leds(2);
    led(3) <= rx_overflow_led   when nios_gpio.led_mode = '0' else not nios_gpio.leds(3);

    -- DAC SPI (data latched on falling edge)
    dac_sclk <= not nios_sclk when nios_gpio.spi_mux = '0' else '0';
    dac_sdi  <= nios_sdio     when nios_gpio.spi_mux = '0' else '0';
    dac_csn  <= nios_ss_n(0)  when nios_gpio.spi_mux = '0' else '1';

    -- ADF SPI (data latched on rising edge)
    adf_sclk <= nios_sclk    when nios_gpio.spi_mux = '1' else '0';
    adf_sdi  <= nios_sdio    when nios_gpio.spi_mux = '1' else '0';
    adf_csn  <= nios_ss_n(1) when nios_gpio.spi_mux = '1' else '1';
    adf_ce   <= nios_gpio.spi_mux;

    nios_sdo <= adf_muxout when ((nios_ss_n(1) = '0') and (nios_gpio.spi_mux = '1'))
                else '0';

    -- Power monitor I2C
    pwr_scl     <= i2c_scl_out when i2c_scl_oen = '0' else 'Z';
    pwr_sda     <= i2c_sda_out when i2c_sda_oen = '0' else 'Z';

    i2c_scl_in  <= pwr_scl;
    i2c_sda_in  <= pwr_sda;

    -- Power mux control
    psu_ctl_d   <= "ZZ";

    -- Expansion clock request/enable
    exp_clock_en <= exp_present and exp_clock_req;

    -- Expansion I2C
    exp_i2c_scl <= 'Z';
    exp_i2c_sda <= 'Z';

    -- Expansion GPIO outputs
    generate_xb_gpio_out : for i in exp_gpio'range generate
        exp_gpio(i) <= nios_xb_gpio_out(i) when nios_xb_gpio_oe(i) = '1' else 'Z';
    end generate;









    -- TX sample fifo
    tx_sample_fifo.aclr   <= tx_reset;
    tx_sample_fifo.wclock <= fx3_pclk_pll;
    tx_sample_fifo.rclock <= tx_clock;
    U_tx_sample_fifo : entity work.tx_fifo
        port map (
            aclr                => tx_sample_fifo.aclr,

            wrclk               => tx_sample_fifo.wclock,
            wrreq               => tx_sample_fifo.wreq,
            data                => tx_sample_fifo.wdata,
            wrempty             => tx_sample_fifo.wempty,
            wrfull              => tx_sample_fifo.wfull,
            wrusedw             => tx_sample_fifo.wused,

            rdclk               => tx_sample_fifo.rclock,
            rdreq               => tx_sample_fifo.rreq,
            q                   => tx_sample_fifo.rdata,
            --rdempty             => tx_sample_fifo.rempty,
            rdempty             => tx_sample_fifo_rempty_untriggered,
            rdfull              => tx_sample_fifo.rfull,
            rdusedw             => tx_sample_fifo.rused
        );

    tx_channel_mux : process( all )
        variable ch     : integer range 0 to 1 := 0;
        variable fifo_i : std_logic_vector(11 downto 0) := (others => '0');
        variable fifo_q : std_logic_vector(11 downto 0) := (others => '0');
        variable valid  : std_logic := '0';
    begin
        if( rising_edge(tx_clock) ) then
            if( channel_sel = '0' ) then
                ch := 0;
            else
                ch := 1;
            end if;

            if( tx_sample_fifo.rempty = '0' ) then
                tx_sample_fifo.rreq <= ad9361.ch(ch).dac.i.valid;
                fifo_i := tx_sample_fifo.rdata(11 downto 0);
                fifo_q := tx_sample_fifo.rdata(27 downto 16);
                valid  := ad9361.ch(ch).dac.i.valid;
            else
                tx_sample_fifo.rreq <= '0';
                fifo_i := (others => '0');
                fifo_q := (others => '0');
                valid  := '0';
            end if;

            ad9361.ch(ch).dac.i.data <= fifo_i & "0000";
            ad9361.ch(ch).dac.q.data <= fifo_q & "0000";

            tx_sample_i     <= resize(signed(fifo_i), tx_sample_i'length);
            tx_sample_q     <= resize(signed(fifo_q), tx_sample_q'length);
            tx_sample_valid <= valid;
        end if;
    end process;

    -- TX meta fifo
    tx_meta_fifo.aclr   <= tx_reset;
    tx_meta_fifo.wclock <= fx3_pclk_pll;
    tx_meta_fifo.rclock <= tx_clock;
    U_tx_meta_fifo : entity work.tx_meta_fifo
        port map (
            aclr                => tx_meta_fifo.aclr,

            wrclk               => tx_meta_fifo.wclock,
            wrreq               => tx_meta_fifo.wreq,
            data                => tx_meta_fifo.wdata,
            wrempty             => tx_meta_fifo.wempty,
            wrfull              => tx_meta_fifo.wfull,
            wrusedw             => tx_meta_fifo.wused,

            rdclk               => tx_meta_fifo.rclock,
            rdreq               => tx_meta_fifo.rreq,
            q                   => tx_meta_fifo.rdata,
            rdempty             => tx_meta_fifo.rempty,
            rdfull              => tx_meta_fifo.rfull,
            rdusedw             => tx_meta_fifo.rused
        );

    --U_fifo_reader : entity work.fifo_reader
    --  port map (
    --    clock               =>  tx_clock,
    --    reset               =>  tx_reset,
    --    enable              =>  tx_enable,
    --
    --    usb_speed           =>  usb_speed_tx,
    --    meta_en             =>  meta_en_tx,
    --    timestamp           =>  tx_timestamp,
    --
    --    fifo_empty          =>  tx_sample_fifo.rempty,
    --    fifo_usedw          =>  tx_sample_fifo.rused,
    --    fifo_data           =>  tx_sample_fifo.rdata,
    --    fifo_read           =>  tx_sample_fifo.rreq,
    --
    --    meta_fifo_empty     =>  tx_meta_fifo.rempty,
    --    meta_fifo_usedw     =>  tx_meta_fifo.rused,
    --    meta_fifo_data      =>  tx_meta_fifo.rdata,
    --    meta_fifo_read      =>  tx_meta_fifo.rreq,
    --
    --    out_i               =>  tx_sample_i,
    --    out_q               =>  tx_sample_q,
    --    out_valid           =>  tx_sample_valid,
    --
    --    underflow_led       =>  tx_underflow_led,
    --    underflow_count     =>  open,
    --    underflow_duration  =>  x"ffff"
    --  ) ;












    -- RX sample fifo
    rx_sample_fifo.aclr   <= not rx_enable_pclk;
    rx_sample_fifo.wclock <= rx_clock;
    rx_sample_fifo.rclock <= fx3_pclk_pll;
    U_rx_sample_fifo : entity work.rx_fifo
        port map (
            aclr                => rx_sample_fifo.aclr,

            wrclk               => rx_sample_fifo.wclock,
            wrreq               => rx_sample_fifo.wreq,
            data                => rx_sample_fifo.wdata,
            wrempty             => rx_sample_fifo.wempty,
            wrfull              => rx_sample_fifo.wfull,
            wrusedw             => rx_sample_fifo.wused,

            rdclk               => rx_sample_fifo.rclock,
            rdreq               => rx_sample_fifo.rreq,
            q                   => rx_sample_fifo.rdata,
            rdempty             => rx_sample_fifo.rempty,
            rdfull              => rx_sample_fifo.rfull,
            rdusedw             => rx_sample_fifo.rused
        );

    -- RX meta fifo
    rx_meta_fifo.aclr   <= not rx_enable_pclk;
    rx_meta_fifo.wclock <= rx_clock;
    rx_meta_fifo.rclock <= fx3_pclk_pll;
    U_rx_meta_fifo : entity work.rx_meta_fifo
        port map (
            aclr                => rx_meta_fifo.aclr,

            wrclk               => rx_meta_fifo.wclock,
            wrreq               => rx_meta_fifo.wreq,
            data                => rx_meta_fifo.wdata,
            wrempty             => rx_meta_fifo.wempty,
            wrfull              => rx_meta_fifo.wfull,
            wrusedw             => rx_meta_fifo.wused,

            rdclk               => rx_meta_fifo.rclock,
            rdreq               => rx_meta_fifo.rreq,
            q                   => rx_meta_fifo.rdata,
            rdempty             => rx_meta_fifo.rempty,
            rdfull              => rx_meta_fifo.rfull,
            rdusedw             => rx_meta_fifo.rused
        );


    -- RX loopback fifo
    rx_loopback_fifo.aclr   <= '1' when tx_reset = '1' or tx_loopback_enabled = '0' else '0';
    rx_loopback_fifo.wclock <= tx_clock;
    rx_loopback_fifo.wdata  <= std_logic_vector(tx_sample_i & tx_sample_q) when tx_loopback_enabled = '1' else (others => '0');
    rx_loopback_fifo.wreq   <= tx_sample_valid when tx_loopback_enabled = '1' else '0';
    rx_loopback_fifo.rclock <= rx_clock;

    U_rx_loopback_fifo : entity work.rx_fifo
        port map (
            aclr                => rx_loopback_fifo.aclr,

            wrclk               => rx_loopback_fifo.wclock,
            wrreq               => rx_loopback_fifo.wreq,
            data                => rx_loopback_fifo.wdata,
            wrempty             => rx_loopback_fifo.wempty,
            wrfull              => rx_loopback_fifo.wfull,
            wrusedw             => rx_loopback_fifo.wused,

            rdclk               => rx_loopback_fifo.rclock,
            rdreq               => rx_loopback_fifo.rreq,
            q                   => rx_loopback_fifo.rdata,
            rdempty             => rx_loopback_fifo.rempty,
            rdfull              => rx_loopback_fifo.rfull,
            rdusedw             => rx_loopback_fifo.rused
        );

    rx_loopback_fifo_out : process( rx_reset, rx_loopback_fifo.rclock )
        constant WATERLINE          : natural := 16;
        variable already_strobed    : boolean := false;
    begin
        if (rx_reset = '1') then
            rx_loopback_enabled     <= '0';
            rx_loopback_fifo.rreq   <= '0';
            rx_loopback_i           <= (others => '0');
            rx_loopback_q           <= (others => '0');
            rx_loopback_valid       <= '0';
        elsif( rising_edge(rx_loopback_fifo.rclock) ) then
            rx_loopback_enabled     <= '0';
            rx_loopback_fifo.rreq   <= '0';
            rx_loopback_i           <= rx_loopback_i;
            rx_loopback_q           <= rx_loopback_q;
            rx_loopback_valid       <= '0';

            -- is loopback enabled?
            if (rx_mux_mode = RX_MUX_DIGITAL_LOOPBACK) then
                rx_loopback_enabled <= rx_enable;
            end if;

            -- do the loopback
            if (rx_loopback_enabled = '1') then
                rx_loopback_i       <= resize(signed(rx_loopback_fifo.rdata(31 downto 16)), rx_loopback_i'length);
                rx_loopback_q       <= resize(signed(rx_loopback_fifo.rdata(15 downto 0)), rx_loopback_q'length);
                rx_loopback_valid   <= rx_loopback_fifo.rreq;
            end if;

            -- read from the fifo if req'd
            if (unsigned(rx_loopback_fifo.rused) > WATERLINE) then
                rx_loopback_fifo.rreq   <= rx_loopback_enabled and not rx_loopback_fifo.rempty;
            end if;

            -- handle situation where fifo is empty but we tried to rreq from it
            if (rx_loopback_fifo.rreq = '1' and already_strobed) then
                already_strobed     := false;
                rx_loopback_valid   <= '0';
            end if;

            -- detect above condition
            already_strobed := (rx_loopback_fifo.rreq = '1' and rx_loopback_fifo.rempty = '1');
        end if;
    end process;










    -- Sample bridges
    U_fifo_writer : entity work.fifo_writer
      port map (
        clock               =>  rx_clock,
        reset               =>  rx_reset,
        enable              =>  rx_enable,

        usb_speed           =>  usb_speed_rx,
        meta_en             =>  meta_en_rx,
        timestamp           =>  rx_timestamp,

        fifo_full           =>  rx_sample_fifo.wfull,
        fifo_usedw          =>  rx_sample_fifo.wused,
        fifo_data           =>  rx_sample_fifo.wdata,
        fifo_write          =>  rx_sample_fifo.wreq,

        meta_fifo_full      =>  rx_meta_fifo.wfull,
        meta_fifo_usedw     =>  rx_meta_fifo.wused,
        meta_fifo_data      =>  rx_meta_fifo.wdata,
        meta_fifo_write     =>  rx_meta_fifo.wreq,

        in_i                =>  resize(rx_mux_i,16),
        in_q                =>  resize(rx_mux_q,16),
        in_valid            =>  rx_mux_valid,

        overflow_led        =>  rx_overflow_led,
        overflow_count      =>  open,
        overflow_duration   =>  x"ffff"
      );

    lms_rx_enable_sig <= rx_enable;

    -- RX Trigger
    rxtrig : entity work.trigger(async)
      generic map (
        DEFAULT_OUTPUT  => '0'
      ) port map (
        armed           => rx_trigger_arm,
        fired           => rx_trigger_fire,
        master          => rx_trigger_master,
        trigger_in      => rx_trigger_line,
        trigger_out     => rx_trigger_line,
        signal_in       => lms_rx_enable_sig,
        signal_out      => rx_trigger_signal_out
      );

    rx_trigger_arm_rb    <= rx_trigger_arm;
    rx_trigger_fire_rb   <= rx_trigger_fire;
    rx_trigger_master_rb <= rx_trigger_master;
    rx_trigger_line_rb   <= rx_trigger_line;
    rx_trigger_unused_rb <= (others => '0');


    txtrig : entity work.trigger(async)
      generic map (
        DEFAULT_OUTPUT  => '1'
      ) port map (
        armed           => tx_trigger_arm_sync,
        fired           => tx_trigger_fire,
        master          => tx_trigger_master,
        trigger_in      => tx_trigger_line_sync,
        trigger_out     => tx_trigger_line,
        signal_in       => tx_sample_fifo_rempty_untriggered,
        signal_out      => tx_sample_fifo.rempty
      );

    tx_trigger_arm_rb    <= tx_trigger_arm;
    tx_trigger_fire_rb   <= tx_trigger_fire;
    tx_trigger_master_rb <= tx_trigger_master;
    tx_trigger_line_rb   <= tx_trigger_line;
    tx_trigger_unused_rb <= (others => '0');


    rx_channel_mux : process( all )
        variable ch : integer range 0 to 1 := 0;
    begin
        if( rising_edge(rx_clock) ) then
            if( channel_sel = '0' ) then
                ch := 0;
            else
                ch := 1;
            end if;

            rx_sample_i(15 downto 12) <= ( others => ad9361.ch(ch).adc.i.data(11) );
            rx_sample_i(11 downto 0)  <= signed(ad9361.ch(ch).adc.i.data(11 downto 0));
            rx_sample_q(15 downto 12) <= ( others => ad9361.ch(ch).adc.q.data(11) );
            rx_sample_q(11 downto 0)  <= signed(ad9361.ch(ch).adc.q.data(11 downto 0));
            rx_sample_valid           <= ad9361.ch(ch).adc.i.valid and
                                         ad9361.ch(ch).adc.q.valid;
        end if;
    end process;


    U_rx_siggen : entity work.signal_generator
      port map (
        clock           =>  rx_clock,
        reset           =>  rx_reset,
        enable          =>  rx_enable,

        mode            =>  rx_gen_mode,

        sample_i        =>  rx_gen_i,
        sample_q        =>  rx_gen_q,
        sample_valid    =>  rx_gen_valid
      );

    rx_mux_mode <= rx_mux_mode_t'val(to_integer(rx_mux_sel));

    rx_mux : process(rx_reset, rx_clock)
    begin
        if( rx_reset = '1' ) then
            rx_mux_i     <= (others =>'0');
            rx_mux_q     <= (others =>'0');
            rx_mux_valid <= '0';
            rx_gen_mode  <= '0';
        elsif( rising_edge(rx_clock) ) then
            case rx_mux_mode is
                when RX_MUX_NORMAL =>
                    rx_mux_i <= rx_sample_i;
                    rx_mux_q <= rx_sample_q;
                    if( lms_rx_enable_qualified = '1' ) then
                        rx_mux_valid <= rx_sample_valid;
                    else
                        rx_mux_valid <= '0';
                    end if;
                when RX_MUX_12BIT_COUNTER | RX_MUX_32BIT_COUNTER =>
                    rx_mux_i     <= rx_gen_i;
                    rx_mux_q     <= rx_gen_q;
                    rx_mux_valid <= rx_gen_valid;
                    if( rx_mux_mode = RX_MUX_32BIT_COUNTER ) then
                        rx_gen_mode <= '1';
                    else
                        rx_gen_mode <= '0';
                    end if;
                when RX_MUX_ENTROPY =>
                    -- Not yet implemented
                    rx_mux_i     <= (others => '0');
                    rx_mux_q     <= (others => '0');
                    rx_mux_valid <= '0';
                when RX_MUX_DIGITAL_LOOPBACK =>
                    rx_mux_i     <= rx_loopback_i;
                    rx_mux_q     <= rx_loopback_q;
                    rx_mux_valid <= rx_loopback_valid;
                when others =>
                    rx_mux_i     <= (others =>'0');
                    rx_mux_q     <= (others =>'0');
                    rx_mux_valid <= '0';
            end case;
        end if;
    end process;







    set_tx_ts_reset : process(tx_clock, tx_reset)
    begin
        if( tx_reset = '1' ) then
            tx_ts_reset <= '1';
        elsif( rising_edge(tx_clock) ) then
            if( meta_en_tx = '1' ) then
                tx_ts_reset <= '0';
            else
                tx_ts_reset <= '1';
            end if;
        end if;
    end process;

    set_rx_ts_reset : process(rx_clock, rx_reset)
    begin
        if( rx_reset = '1' ) then
            rx_ts_reset <= '1';
        elsif( rising_edge(rx_clock) ) then
            if( meta_en_rx = '1' ) then
                rx_ts_reset <= '0';
            else
                rx_ts_reset <= '1';
            end if;
        end if;
    end process;


    -- ========================================================================
    -- RESET SYNCHRONIZERS
    -- ========================================================================

    U_reset_sync_pclk : entity work.reset_synchronizer
        generic map (
            INPUT_LEVEL         =>  '1',
            OUTPUT_LEVEL        =>  '1'
        )
        port map (
            clock               =>  fx3_pclk_pll,
            async               =>  sys_reset_async,
            sync                =>  sys_reset_pclk
        );

    U_reset_sync_sys : entity work.reset_synchronizer
        generic map (
            INPUT_LEVEL         =>  '1',
            OUTPUT_LEVEL        =>  '1'
        )
        port map (
            clock               =>  sys_clock,
            async               =>  sys_reset_async,
            sync                =>  sys_reset
        );

    U_reset_sync_rx : entity work.reset_synchronizer
        generic map (
            INPUT_LEVEL         =>  '1',
            OUTPUT_LEVEL        =>  '1'
        )
        port map (
            clock               =>  rx_clock,
            async               =>  sys_reset_pclk,
            sync                =>  rx_reset
        );

    U_reset_sync_tx : entity work.reset_synchronizer
        generic map (
            INPUT_LEVEL         =>  '1',
            OUTPUT_LEVEL        =>  '1'
        )
        port map (
            clock               =>  tx_clock,
            async               =>  sys_reset_pclk,
            sync                =>  tx_reset
        );

    U_reset_sync_loopback : entity work.reset_synchronizer
        generic map (
            INPUT_LEVEL         => '0',
            OUTPUT_LEVEL        => '0'
        )
        port map (
            clock               =>  tx_clock,
            async               =>  rx_loopback_enabled,
            sync                =>  tx_loopback_enabled
        );

    U_reset_sync_tx_trig_arm : entity work.reset_synchronizer
        generic map (
            INPUT_LEVEL     =>  '0',
            OUTPUT_LEVEL    =>  '0'
        )
        port map (
            clock           =>  tx_clock,
            async           =>  tx_trigger_arm,
            sync            =>  tx_trigger_arm_sync
        );


    -- ========================================================================
    -- SYNCHRONIZERS
    -- ========================================================================

    U_sync_usb_speed_pclk : entity work.synchronizer
        generic map (
            RESET_LEVEL         =>  '0'
        )
        port map (
            reset               =>  '0',
            clock               =>  fx3_pclk_pll,
            async               =>  nios_gpio.usb_speed,
            sync                =>  usb_speed_pclk
        );

    U_sync_usb_speed_rx : entity work.synchronizer
        generic map (
            RESET_LEVEL         =>  '0'
        )
        port map (
            reset               =>  '0',
            clock               =>  rx_clock,
            async               =>  nios_gpio.usb_speed,
            sync                =>  usb_speed_rx
        );

    U_sync_usb_speed_tx : entity work.synchronizer
        generic map (
            RESET_LEVEL         =>  '0'
        )
        port map (
            reset               =>  '0',
            clock               =>  tx_clock,
            async               =>  nios_gpio.usb_speed,
            sync                =>  usb_speed_tx
        );


    U_sync_meta_en_pclk : entity work.synchronizer
        generic map (
            RESET_LEVEL         =>  '0'
        )
        port map (
            reset               =>  '0',
            clock               =>  fx3_pclk_pll,
            async               =>  nios_gpio.meta_sync,
            sync                =>  meta_en_pclk
        );

    U_sync_meta_en_rx : entity work.synchronizer
        generic map (
            RESET_LEVEL         =>  '0'
        )
        port map (
            reset               =>  '0',
            clock               =>  rx_clock,
            async               =>  nios_gpio.meta_sync,
            sync                =>  meta_en_rx
        );

    U_sync_meta_en_tx : entity work.synchronizer
        generic map (
            RESET_LEVEL         =>  '0'
        )
        port map (
            reset               =>  '0',
            clock               =>  tx_clock,
            async               =>  nios_gpio.meta_sync,
            sync                =>  meta_en_tx
        );

    generate_sync_rx_mux_sel : for i in rx_mux_sel'range generate
        U_sync_rx_mux_sel : entity work.synchronizer
            generic map (
                RESET_LEVEL         =>  '0'
            )
            port map (
                reset               =>  '0',
                clock               =>  rx_clock,
                async               =>  nios_gpio.rx_mux_sel(i),
                sync                =>  rx_mux_sel(i)
            );
    end generate;

    U_sync_channel_sel : entity work.synchronizer
        generic map (
            RESET_LEVEL         =>  '0'
        )
        port map (
            reset               =>  '0',
            clock               =>  rx_clock,
            async               =>  nios_gpio.channel_sel,
            sync                =>  channel_sel
        );

    generate_sync_adi_ctrl_out : for i in adi_ctrl_out'range generate
        U_sync_adi_ctrl_out : entity work.synchronizer
            generic map (
                RESET_LEVEL         =>  '0'
            )
            port map (
                reset               =>  '0',
                clock               =>  sys_clock,
                async               =>  adi_ctrl_out(i),
                sync                =>  rffe_gpio.i.ctrl_out(i)
            );
    end generate;

    generate_sync_xb_gpio_in : for i in exp_gpio'range generate
        U_sync_xb_gpio_in : entity work.synchronizer
          generic map (
            RESET_LEVEL         =>  '0'
          ) port map (
            reset               =>  '0',
            clock               =>  sys_clock,
            async               =>  exp_gpio(i),
            sync                =>  nios_xb_gpio_in(i)
          );
    end generate;

    U_sync_rx_enable : entity work.synchronizer
        generic map (
            RESET_LEVEL =>  '0'
        )
        port map (
            reset       =>  rx_reset,
            clock       =>  rx_clock,
            async       =>  rx_enable_pclk,
            sync        =>  rx_enable
        );

    U_sync_tx_enable : entity work.synchronizer
        generic map (
            RESET_LEVEL =>  '0'
        )
        port map (
            reset       =>  tx_reset,
            clock       =>  tx_clock,
            async       =>  tx_enable_pclk,
            sync        =>  tx_enable
        );

    U_sync_rx_trig_signal_out : entity work.synchronizer
        generic map (
            RESET_LEVEL =>  '0'
        )
        port map (
            reset       =>  rx_reset,
            clock       =>  rx_clock,
            async       =>  rx_trigger_signal_out,
            sync        =>  lms_rx_enable_qualified
        );

    U_sync_tx_trig_trigger_line : entity work.synchronizer
        generic map (
            RESET_LEVEL =>  '0'
        )
        port map (
            reset       =>  tx_reset,
            clock       =>  tx_clock,
            async       =>  tx_trigger_line,
            sync        =>  tx_trigger_line_sync
        );


    -- ========================================================================
    -- HANDSHAKES
    -- ========================================================================

    drive_handshake_timestamp : process( fx3_pclk_pll, sys_reset_pclk )
    begin
        if( sys_reset_pclk = '1' ) then
            timestamp_req <= '0';
        elsif( rising_edge(fx3_pclk_pll) ) then
            if( meta_en_pclk = '0' ) then
                timestamp_req <= '0';
            else
                if( timestamp_ack = '0' ) then
                    timestamp_req <= '1';
                elsif( timestamp_ack = '1' ) then
                    timestamp_req <= '0';
                end if;
            end if;
        end if;
    end process;

    U_handshake_timestamp : entity work.handshake
        generic map (
            DATA_WIDTH          =>  tx_timestamp'length
        )
        port map (
            source_clock        =>  tx_clock,
            source_reset        =>  tx_reset,
            source_data         =>  std_logic_vector(tx_timestamp),

            dest_clock          =>  fx3_pclk_pll,
            dest_reset          =>  sys_reset_pclk,
            unsigned(dest_data) =>  fx3_timestamp,
            dest_req            =>  timestamp_req,
            dest_ack            =>  timestamp_ack
        );

end architecture;
